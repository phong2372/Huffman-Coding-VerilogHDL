`timescale 1ns/1ps
module huffman_test;

	// Inputs
	reg CLK;
	reg nRST;
	reg [3:0] in;
	reg start;

	// Outputs
	wire done;
	wire	[10:0] length;

	huffman dut(
	.CLK(CLK),
	.nRST(nRST),
	.start(start),
	.in(in),
	.length(length),
	.done(done)
	);
	
	//integer K;

	initial begin
		// Initialize Inputs
		CLK = 0;
		nRST = 0;
		in = 4'b0000;
		//in <= 1024'b0101_0101_0101_0100_0101_0100_0101_0100_0011_0101_0100_0011_0010_0101_0100_0011_0010_0101_0100_0011_0010_0101_0100_0011_0010_0001_0101_0100_0011_0010_0001;
		//in <= 1024'b1010_1010_1010_1001_1010_1001_1010_1001_1000_1010_1001_1000_1010_1001_1000_0111_1010_1001_1000_0111_1010_1001_1000_0111_0110_1010_1001_1000_0111_0110_1010_1001_1000_0111_0110_0101_1010_1001_1000_0111_0110_0101_1010_1001_1000_0111_0110_0101_0100_1010_1001_1000_0111_0110_0101_0100_1010_1001_1000_0111_0110_0101_0100_0011_1010_1001_1000_0111_0110_0101_0100_0011_1010_1001_1000_0111_0110_0101_0100_0011_0010_1010_1001_1000_0111_0110_0101_0100_0011_0010_1010_1001_1000_0111_0110_0101_0100_0011_0010_0001_1010_1001_1000_0111_0110_0101_0100_0011_0010_0001_1010_1001_1000_0111_0110_0101_0100_0011_0010_0001_1010_1010_1010_1001_1010_1001_1010_1001_1000_1010_1001_1000_1010_1001_1000_0111_1010_1001_1000_0111_1010_1001_1000_0111_0110_1010_1001_1000_0111_0110_1010_1001_1000_0111_0110_0101_1010_1001_1000_0111_0110_0101_1010_1001_1000_0111_0110_0101_0100_1010_1001_1000_0111_0110_0101_0100_1010_1001_1000_0111_0110_0101_0100_0011_1010_1001_1000_0111_0110_0101_0100_0011_1010_1001_1000_0111_0110_0101_0100_0011_0010_1010_1001_1000_0111_0110_0101_0100_0011_0010_1010_1001_1000_0111_0110_0101_0100_0011_0010_0001_1010_1001_1000_0111_0110_0101_0100_0011_0010_0001_1010_1001_1000_0111_0110_0101_0100_0011_0010_0001;

		// Wait 100 ns for global reset to finish
		#100;      
		nRST = 1;
		#5;
		start = 1;
 	end
	parameter DELAY = 1;
	always 
		#DELAY CLK = ~ CLK;
	

endmodule

